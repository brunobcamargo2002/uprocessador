library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
    port(
        clk: in std_logic;
        address: in unsigned(6 downto 0);
        data: out unsigned(15 downto 0)
    );
end entity;




architecture a_rom of rom is
    type mem is array(0 to 127) of unsigned(15 downto 0);
    constant content: mem :=(
        1 => B"0001_001_000000000", -- ld r1, 0
        2 => B"0001_010_000100000", -- ld r2, 32
        3 => B"0110_000_001_000000", -- mova r1
        4 => B"0011_000_000000001", -- addi 1
        5 => B"0111_001_000000000", -- movr r1
        6 => B"1101_000_001_000000", -- sw r1
        7 => B"0110_000_001_000000", -- mova r1
        8 => B"0100_000_010_000000", -- sub r2
        9 => B"1011_1111010_00000", -- jc -6
-----------------------------------------------------
-------------Crivo de Eratóstenes -------------------
-----------------------------------------------------
        10 => B"0001_001_000000010", -- ld r1, 2
        11 => B"0001_010_000100000", -- ld r2, 32
        12 => B"0110_000_001_000000", -- mova r1
        13 => B"0011_000_000000010", -- addi 2
        14 => B"0111_001_000000000", -- movr r1
        15 => B"1101_000_000_000000", -- sw r0
        16 => B"0110_000_001_000000", -- mova r1
        17 => B"0100_000_010_000000", -- sub r2
        18 => B"1011_1111010_00000", -- jc -6

        19 => B"0001_001_000000001", -- ld r1, 1
        20 => B"0110_000_000_000000", -- mova r0
        21 => B"0010_000_001_000000", -- add r1
        22 => B"0011_000_000000010", -- addi 2
        23 => B"0111_001_000000000", -- movr r1
        24 => B"1100_011_000000000", -- lw r3 --
        25 => B"0110_000_011_000000", -- mova r3
        26 => B"1001_1111010_00000", -- jz -6
        


        27 => B"0110_000_001_000000", -- mova r1
        28 => B"0010_000_001_000000", -- add r1
        29 => B"0010_000_001_000000", -- add r1
        30 => B"0111_011_000000000", -- movr r3
        31 => B"0110_000_011_000000", -- mova r3
        32 => B"1101_000_000_000000", -- sw r0
        33 => B"0010_000_001_000000", -- add r1
        34 => B"0010_000_001_000000", -- add r1
        35 => B"0111_011_000000000", -- movr r3
        36 => B"0100_000_010_000000", -- sub r2
        37 => B"1011_1111010_00000", -- jc -6

        38 => B"0110_000_001_000000", -- mova r1
        39 => B"0011_000_000000010", -- addi 2
        40 => B"0111_001_000000000", -- movr r1
        41 => B"0100_000_010_000000", -- sub r2
        42 => B"1011_1101110_00000", -- jc -18

        43 => B"0001_100_000000000", -- ld r4, 0
        44 => B"0110_000_100_000000", -- mova r4
        45 => B"0011_000_000000001", -- addi, 1
        46 => B"1100_101_000000000", -- lw r5
        47 => B"0111_100_000000000", -- movr r4
        48 => B"0100_000_010_000000", -- sub r2
        49 => B"1011_1111011_00000", -- jc -5

        others => (others=>'0')
    );
begin
    process(clk)
    begin
        if(rising_edge(clk)) then
            data <= content(to_integer(address));
        end if;
    end process;
end architecture;
