library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
    port(
        clk: in std_logic;
        address: in unsigned(6 downto 0);
        data: out unsigned(15 downto 0)
    );
end entity;




architecture a_rom of rom is
    type mem is array(0 to 127) of unsigned(15 downto 0);
    constant content: mem :=(
        -- Carregar 19563_10 = 4C6B_16 em r4 --
        1 => B"0001_001_000000000", -- ld r1, 0 -- iterador
        2 => B"0001_010_100000000", -- ld r2, 256 -- op mult 1
        3 => B"0001_011_001001110", -- ld r3, 78 -- op mult 2
        4 => B"0001_100_000000000", -- ld r4, 0 -- resultado
        5 => B"0110_000_100_000000", -- mova r4
        6 => B"0010_000_010_000000", -- add r2
        7 => B"0111_100_0000_00000", -- mvr r4
        8 => B"0110_000_001_000000", -- mova r1
        9 => B"0011_000_000000001", -- addi 1
        10 => B"1110_000_011_000000", -- cmp r3
        11 => B"0111_001_0000_00000", -- mvr r1
        12 => B"1011_1111001_00000", -- jc -7
        13 => B"0110_000_100_000000", -- mova r4
        -- 14 => B"0101_000_00000_0001", -- subi 1
        14 => B"0111_010_0000_00000", -- mvr r2
        15 => B"0001_100_000000000", -- ld r4, 0
        16 => B"0001_011_000000000", -- ld r3, 0

        17 => B"0001_001_000000000", -- ld r1, 0
        18 => B"0110_000_001_000000", -- mova r1
        19 => B"0011_000_000000001", -- addi 1
        20 => B"0111_001_000000000", -- movr r1
        21 => B"1101_000_001_000000", -- sw r1
        22 => B"0110_000_001_000000", -- mova r1
        23 => B"0100_000_010_000000", -- sub r2
        24 => B"1011_1111010_00000", -- jc -6
-----------------------------------------------------
-------------Crivo de Eratóstenes -------------------
-----------------------------------------------------
-- Remove os pares (eu acho) --
        25 => B"0001_001_000000010", -- ld r1, 2
        26 => B"0110_000_001_000000", -- mova r1
        27 => B"0011_000_000000010", -- addi 2
        28 => B"0111_001_000000000", -- movr r1
        29 => B"1101_000_000_000000", -- sw r0
        30 => B"0110_000_001_000000", -- mova r1
        31 => B"0100_000_010_000000", -- sub r2
        32 => B"1011_1111010_00000", -- jc -6


        33 => B"0001_001_000000001", -- ld r1, 1
        34 => B"0110_000_000_000000", -- mova r0
        35 => B"0010_000_001_000000", -- add r1
        36 => B"0011_000_000000010", -- addi 2
        37 => B"0111_001_000000000", -- movr r1
        38 => B"1100_011_000000000", -- lw r3 --
        39 => B"0110_000_011_000000", -- mova r3
        40 => B"1001_1111010_00000", -- jz -6
       


        41 => B"0110_000_001_000000", -- mova r1
        42 => B"0010_000_001_000000", -- add r1
        43 => B"0010_000_001_000000", -- add r1
        44 => B"0111_011_000000000", -- movr r3
        45 => B"0110_000_011_000000", -- mova r3
        46 => B"1101_000_000_000000", -- sw r0
        47 => B"0010_000_001_000000", -- add r1
        48 => B"0010_000_001_000000", -- add r1
        49 => B"0111_011_000000000", -- movr r3
        50 => B"0100_000_010_000000", -- sub r2
        51 => B"1011_1111010_00000", -- jc -6

        52 => B"0110_000_001_000000", -- mova r1
        53 => B"0011_000_000000010", -- addi 2
        54 => B"0111_001_000000000", -- movr r1
        55 => B"0100_000_010_000000", -- sub r2
        56 => B"1011_1101110_00000", -- jc -18

        57 => B"0001_100_000000000", -- ld r4, 0
        58 => B"0110_000_100_000000", -- mova r4
        59 => B"0011_000_000000001", -- addi, 1
        60 => B"1100_101_000000000", -- lw r5
        61 => B"0111_100_000000000", -- movr r4
        62 => B"0100_000_010_000000", -- sub r2
        63 => B"1011_1111011_00000", -- jc -5

        others => (others=>'0')
    );
begin
    process(clk)
    begin
        if(rising_edge(clk)) then
            data <= content(to_integer(address));
        end if;
    end process;
end architecture;
